module hello
  (input clk_i
  ,input reset_i);

   initial 
     $display("Hello World!");

endmodule
